`ifndef _inst_mem_v_
`define _inst_mem_v_
`endif

module inst_mem(addr, data);
  input wire [31:0] addr;
  output reg [31:0] data;

  reg [31:0] rf_data [127:0];

  always @(addr)
    data = rf_data[addr[6:0]];
    
  // lab 1 instruction memory data test
  /*
  initial begin
    rf_data[0] <= 32'hA00000AA;
    rf_data[1] <= 32'h10000011;
    rf_data[2] <= 32'h20000022;
    rf_data[3] <= 32'h30000033;
    rf_data[4] <= 32'h40000044;
    rf_data[5] <= 32'h50000055;
    rf_data[6] <= 32'h60000066;
    rf_data[7] <= 32'h70000077;
    rf_data[8] <= 32'h80000088;
    rf_data[9] <= 32'h90000099;
  end
  */
  
  // lab 2 instruction memory data test
  /*
  initial begin
    rf_data[0] <= 32'h002300aa;
    rf_data[1] <= 32'h10254321;
    rf_data[2] <= 32'h00200022;
    rf_data[3] <= 32'h8c123456;
    rf_data[4] <= 32'h8f123456;
    rf_data[5] <= 32'had654321;
    rf_data[6] <= 32'h13012345;
    rf_data[7] <= 32'hac654321;
    rf_data[8] <= 32'h12012345;
  end
  */
  
  
  // lab 3 instuction memory data test
  /*
  initial begin
    rf_data[0] <= 32'h002300AA;
    rf_data[1] <= 32'h10654321;
    rf_data[2] <= 32'h00100022;
    rf_data[3] <= 32'h8C123456;
    rf_data[4] <= 32'h8F123456;
    rf_data[5] <= 32'hAD654321;
    rf_data[6] <= 32'h13012345;
    rf_data[7] <= 32'hAC654321;
    rf_data[8] <= 32'h12012345;
  end
  */
  
  // lab 4 instruction memory data test
  
  //initial begin
   // rf_data[0] <= 32'h00221820;
   // rf_data[1] <= 32'h8C220004;
   // rf_data[2] <= 32'b101011_00001_00010_00000_00000_000100;
   // rf_data[3] <= 32'h8C220004;
        //rf_data[2] <= 32'hACC50008;
    //rf_data[3] <= 32'h10000000;
    //rf_data[3] <= 32'b000100_00000_00000_11111_11111_111100;
  //end
  
  // instructions for final test
  initial begin
    rf_data[0] = 32'b100011_00000_00001_0000_0000_0000_0001;    //_LW_r_1_,_1(_r0_)
    rf_data[1] = 32'b100011_00000_00010_0000_0000_0000_0010;    //LW_r_2_,_2(_r0_)
    rf_data[2] = 32'b100011_00000_00011_0000_0000_0000_0011;    //LW_r_3_,_3(_r0_)
    rf_data[3] = 32'b1000_0000_0000_0000_0000_0000_0000_0000;    //NOP
    rf_data[4] = 32'b1000_0000_0000_0000_0000_0000_0000_0000;    //NOP
    rf_data[5] = 32'b000000_00001_00010_00001_00000_100000;    //ADD_r_1_,_r_1_,_r2
    rf_data[6] = 32'b1000_0000_0000_0000_0000_0000_0000_0000;    //NOP
    rf_data[7] = 32'b1000_0000_0000_0000_0000_0000_0000_0000;    //NOP
    rf_data[8] = 32'b1000_0000_0000_0000_0000_0000_0000_0000;    //NOP
    rf_data[9] = 32'b000000_00001_00011_00001_00000_100000;    //ADD_r_1_,_r_1_,_r3
    rf_data[10] = 32'b1000_0000_0000_0000_0000_0000_0000_0000;    //NOP
    rf_data[11] = 32'b1000_0000_0000_0000_0000_0000_0000_0000;    //NOP
    rf_data[12] = 32'b1000_0000_0000_0000_0000_0000_0000_0000;    //NOP
    rf_data[13] = 32'b000000_00001_00001_00001_00000_100000;    //ADD_r_1_,_r_1_,_r1
    rf_data[14] = 32'b1000_0000_0000_0000_0000_0000_0000_0000;    //NOP
    rf_data[15] = 32'b1000_0000_0000_0000_0000_0000_0000_0000;    //NOP
    rf_data[16] = 32'b1000_0000_0000_0000_0000_0000_0000_0000;    //NOP
    rf_data[17] = 32'b1000_0000_0000_0000_0000_0000_0000_0000;    //NOP
    rf_data[18] = 32'b000000_00001_00000_00001_00000_100000;    //ADD_r_1_,_r_1_,_r0
    rf_data[19] = 32'b1000_0000_0000_0000_0000_0000_0000_0000;    //NOP
    rf_data[20] = 32'b1000_0000_0000_0000_0000_0000_0000_0000;    //NOP
    rf_data[21] = 32'b1000_0000_0000_0000_0000_0000_0000_0000;    //NOP
    rf_data[22] = 32'b1000_0000_0000_0000_0000_0000_0000_0000;    //NOP
    rf_data[23] = 32'b1000_0000_0000_0000_0000_0000_0000_0000;    //NOP
    rf_data[23] = 32'b1000_0000_0000_0000_0000_0000_0000_0000;    //NOP
    rf_data[24] = 32'b000000_00001_00000_00001_00000_100000;    //ADD_r_1_,_r_1_,_r0
  end
  
  
  
  
endmodule